module torrent

struct Peer {
	ip_addr string
	port    int
}
